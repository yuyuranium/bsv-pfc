../../vendor/bluecheck/BlueCheck.bsv